module PingPong ();

// structure
//
// hdmi_sync
// render
// ball
// paddle
// game_state
//
//
endmodule

